LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY intra16x16_datapath IS
  PORT (
  
  );

END intra16x16_datapath;

ARCHITECTURE Behavioral OF intra16x16_datapath IS

BEGIN

END Behavioral;
    
